package DefaultValue ;

// Default Value package
// This package has been moved to the Prelude

endpackage
