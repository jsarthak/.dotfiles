package Contexts;

import ModuleContext::*;
import ModuleCollect::*;

import CBus::*;
import LBus::*;



export ModuleContext::*;
export ModuleCollect::*;

endpackage
